`define DES
//`define SVA